
module Shifter( dataA, dataB, dataOut );
input [31:0] dataA ;
input [4:0] dataB ; // dataA -> 可能被移位的資料 // dataB -> 移幾位元
output [31:0] dataOut ;
wire [31:0] temp1, temp2, temp3, temp4, temp5 ;

  Mux_1 B0_Mux0( .out( temp1[0] ), .in0( dataA[0] ), .in1( 1'b0 ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux1( .out( temp1[1] ), .in0( dataA[1] ), .in1( dataA[0] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux2( .out( temp1[2] ), .in0( dataA[2] ), .in1( dataA[1] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux3( .out( temp1[3] ), .in0( dataA[3] ), .in1( dataA[2] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux4( .out( temp1[4] ), .in0( dataA[4] ), .in1( dataA[3] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux5( .out( temp1[5] ), .in0( dataA[5] ), .in1( dataA[4] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux6( .out( temp1[6] ), .in0( dataA[6] ), .in1( dataA[5] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux7( .out( temp1[7] ), .in0( dataA[7] ), .in1( dataA[6] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux8( .out( temp1[8] ), .in0( dataA[8] ), .in1( dataA[7] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux9( .out( temp1[9] ), .in0( dataA[9] ), .in1( dataA[8] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux10( .out( temp1[10] ), .in0( dataA[10] ), .in1( dataA[9] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux11( .out( temp1[11] ), .in0( dataA[11] ), .in1( dataA[10] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux12( .out( temp1[12] ), .in0( dataA[12] ), .in1( dataA[11] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux13( .out( temp1[13] ), .in0( dataA[13] ), .in1( dataA[12] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux14( .out( temp1[14] ), .in0( dataA[14] ), .in1( dataA[13] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux15( .out( temp1[15] ), .in0( dataA[15] ), .in1( dataA[14] ), .sel( dataB[0] ) ) ; 
  Mux_1 B0_Mux16( .out( temp1[16] ), .in0( dataA[16] ), .in1( dataA[15] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux17( .out( temp1[17] ), .in0( dataA[17] ), .in1( dataA[16] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux18( .out( temp1[18] ), .in0( dataA[18] ), .in1( dataA[17] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux19( .out( temp1[19] ), .in0( dataA[19] ), .in1( dataA[18] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux20( .out( temp1[20] ), .in0( dataA[20] ), .in1( dataA[19] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux21( .out( temp1[21] ), .in0( dataA[21] ), .in1( dataA[20] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux22( .out( temp1[22] ), .in0( dataA[22] ), .in1( dataA[21] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux23( .out( temp1[23] ), .in0( dataA[23] ), .in1( dataA[22] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux24( .out( temp1[24] ), .in0( dataA[24] ), .in1( dataA[23] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux25( .out( temp1[25] ), .in0( dataA[25] ), .in1( dataA[24] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux26( .out( temp1[26] ), .in0( dataA[26] ), .in1( dataA[25] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux27( .out( temp1[27] ), .in0( dataA[27] ), .in1( dataA[26] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux28( .out( temp1[28] ), .in0( dataA[28] ), .in1( dataA[27] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux29( .out( temp1[29] ), .in0( dataA[29] ), .in1( dataA[28] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux30( .out( temp1[30] ), .in0( dataA[30] ), .in1( dataA[29] ), .sel( dataB[0] ) ) ;
  Mux_1 B0_Mux31( .out( temp1[31] ), .in0( dataA[31] ), .in1( dataA[30] ), .sel( dataB[0] ) ) ;
  
  Mux_1 B1_Mux0( .out( temp2[0] ), .in0( temp1[0] ), .in1( 1'b0 ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux1( .out( temp2[1] ), .in0( temp1[1] ), .in1( 1'b0 ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux2( .out( temp2[2] ), .in0( temp1[2] ), .in1( temp1[0] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux3( .out( temp2[3] ), .in0( temp1[3] ), .in1( temp1[1] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux4( .out( temp2[4] ), .in0( temp1[4] ), .in1( temp1[2] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux5( .out( temp2[5] ), .in0( temp1[5] ), .in1( temp1[3] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux6( .out( temp2[6] ), .in0( temp1[6] ), .in1( temp1[4] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux7( .out( temp2[7] ), .in0( temp1[7] ), .in1( temp1[5] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux8( .out( temp2[8] ), .in0( temp1[8] ), .in1( temp1[6] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux9( .out( temp2[9] ), .in0( temp1[9] ), .in1( temp1[7] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux10( .out( temp2[10] ), .in0( temp1[10] ), .in1( temp1[8] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux11( .out( temp2[11] ), .in0( temp1[11] ), .in1( temp1[9] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux12( .out( temp2[12] ), .in0( temp1[12] ), .in1( temp1[10] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux13( .out( temp2[13] ), .in0( temp1[13] ), .in1( temp1[11] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux14( .out( temp2[14] ), .in0( temp1[14] ), .in1( temp1[12] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux15( .out( temp2[15] ), .in0( temp1[15] ), .in1( temp1[13] ), .sel( dataB[1] ) ) ; 
  Mux_1 B1_Mux16( .out( temp2[16] ), .in0( temp1[16] ), .in1( temp1[14] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux17( .out( temp2[17] ), .in0( temp1[17] ), .in1( temp1[15] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux18( .out( temp2[18] ), .in0( temp1[18] ), .in1( temp1[16] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux19( .out( temp2[19] ), .in0( temp1[19] ), .in1( temp1[17] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux20( .out( temp2[20] ), .in0( temp1[20] ), .in1( temp1[18] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux21( .out( temp2[21] ), .in0( temp1[21] ), .in1( temp1[19] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux22( .out( temp2[22] ), .in0( temp1[22] ), .in1( temp1[10] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux23( .out( temp2[23] ), .in0( temp1[23] ), .in1( temp1[21] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux24( .out( temp2[24] ), .in0( temp1[24] ), .in1( temp1[22] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux25( .out( temp2[25] ), .in0( temp1[25] ), .in1( temp1[23] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux26( .out( temp2[26] ), .in0( temp1[26] ), .in1( temp1[24] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux27( .out( temp2[27] ), .in0( temp1[27] ), .in1( temp1[25] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux28( .out( temp2[28] ), .in0( temp1[28] ), .in1( temp1[26] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux29( .out( temp2[29] ), .in0( temp1[29] ), .in1( temp1[27] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux30( .out( temp2[30] ), .in0( temp1[30] ), .in1( temp1[28] ), .sel( dataB[1] ) ) ;
  Mux_1 B1_Mux31( .out( temp2[31] ), .in0( temp1[31] ), .in1( temp1[29] ), .sel( dataB[1] ) ) ;
  
  Mux_1 B2_Mux0( .out( temp3[0] ), .in0( temp2[0] ), .in1( 1'b0 ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux1( .out( temp3[1] ), .in0( temp2[1] ), .in1( 1'b0 ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux2( .out( temp3[2] ), .in0( temp2[2] ), .in1( 1'b0 ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux3( .out( temp3[3] ), .in0( temp2[3] ), .in1( 1'b0 ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux4( .out( temp3[4] ), .in0( temp2[4] ), .in1( temp2[0] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux5( .out( temp3[5] ), .in0( temp2[5] ), .in1( temp2[1] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux6( .out( temp3[6] ), .in0( temp2[6] ), .in1( temp2[2] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux7( .out( temp3[7] ), .in0( temp2[7] ), .in1( temp2[3] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux8( .out( temp3[8] ), .in0( temp2[8] ), .in1( temp2[4] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux9( .out( temp3[9] ), .in0( temp2[9] ), .in1( temp2[5] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux10( .out( temp3[10] ), .in0( temp2[10] ), .in1( temp2[6] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux11( .out( temp3[11] ), .in0( temp2[11] ), .in1( temp2[7] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux12( .out( temp3[12] ), .in0( temp2[12] ), .in1( temp2[8] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux13( .out( temp3[13] ), .in0( temp2[13] ), .in1( temp2[9] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux14( .out( temp3[14] ), .in0( temp2[14] ), .in1( temp2[10] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux15( .out( temp3[15] ), .in0( temp2[15] ), .in1( temp2[11] ), .sel( dataB[2] ) ) ; 
  Mux_1 B2_Mux16( .out( temp3[16] ), .in0( temp2[16] ), .in1( temp2[12] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux17( .out( temp3[17] ), .in0( temp2[17] ), .in1( temp2[13] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux18( .out( temp3[18] ), .in0( temp2[18] ), .in1( temp2[14] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux19( .out( temp3[19] ), .in0( temp2[19] ), .in1( temp2[15] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux20( .out( temp3[20] ), .in0( temp2[20] ), .in1( temp2[16] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux21( .out( temp3[21] ), .in0( temp2[21] ), .in1( temp2[17] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux22( .out( temp3[22] ), .in0( temp2[22] ), .in1( temp2[18] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux23( .out( temp3[23] ), .in0( temp2[23] ), .in1( temp2[19] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux24( .out( temp3[24] ), .in0( temp2[24] ), .in1( temp2[20] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux25( .out( temp3[25] ), .in0( temp2[25] ), .in1( temp2[21] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux26( .out( temp3[26] ), .in0( temp2[26] ), .in1( temp2[22] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux27( .out( temp3[27] ), .in0( temp2[27] ), .in1( temp2[23] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux28( .out( temp3[28] ), .in0( temp2[28] ), .in1( temp2[24] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux29( .out( temp3[29] ), .in0( temp2[29] ), .in1( temp2[25] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux30( .out( temp3[30] ), .in0( temp2[30] ), .in1( temp2[26] ), .sel( dataB[2] ) ) ;
  Mux_1 B2_Mux31( .out( temp3[31] ), .in0( temp2[31] ), .in1( temp2[27] ), .sel( dataB[2] ) ) ;
  
  Mux_1 B3_Mux0( .out( temp4[0] ), .in0( temp3[0] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux1( .out( temp4[1] ), .in0( temp3[1] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux2( .out( temp4[2] ), .in0( temp3[2] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux3( .out( temp4[3] ), .in0( temp3[3] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux4( .out( temp4[4] ), .in0( temp3[4] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux5( .out( temp4[5] ), .in0( temp3[5] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux6( .out( temp4[6] ), .in0( temp3[6] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux7( .out( temp4[7] ), .in0( temp3[7] ), .in1( 1'b0 ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux8( .out( temp4[8] ), .in0( temp3[8] ), .in1( temp3[0] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux9( .out( temp4[9] ), .in0( temp3[9] ), .in1( temp3[1] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux10( .out( temp4[10] ), .in0( temp3[10] ), .in1( temp3[2] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux11( .out( temp4[11] ), .in0( temp3[11] ), .in1( temp3[3] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux12( .out( temp4[12] ), .in0( temp3[12] ), .in1( temp3[4] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux13( .out( temp4[13] ), .in0( temp3[13] ), .in1( temp3[5] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux14( .out( temp4[14] ), .in0( temp3[14] ), .in1( temp3[6] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux15( .out( temp4[15] ), .in0( temp3[15] ), .in1( temp3[7] ), .sel( dataB[3] ) ) ; 
  Mux_1 B3_Mux16( .out( temp4[16] ), .in0( temp3[16] ), .in1( temp3[8] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux17( .out( temp4[17] ), .in0( temp3[17] ), .in1( temp3[9] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux18( .out( temp4[18] ), .in0( temp3[18] ), .in1( temp3[10] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux19( .out( temp4[19] ), .in0( temp3[19] ), .in1( temp3[11] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux20( .out( temp4[20] ), .in0( temp3[20] ), .in1( temp3[12] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux21( .out( temp4[21] ), .in0( temp3[21] ), .in1( temp3[13] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux22( .out( temp4[22] ), .in0( temp3[22] ), .in1( temp3[14] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux23( .out( temp4[23] ), .in0( temp3[23] ), .in1( temp3[15] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux24( .out( temp4[24] ), .in0( temp3[24] ), .in1( temp3[16] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux25( .out( temp4[25] ), .in0( temp3[25] ), .in1( temp3[17] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux26( .out( temp4[26] ), .in0( temp3[26] ), .in1( temp3[18] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux27( .out( temp4[27] ), .in0( temp3[27] ), .in1( temp3[19] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux28( .out( temp4[28] ), .in0( temp3[28] ), .in1( temp3[20] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux29( .out( temp4[29] ), .in0( temp3[29] ), .in1( temp3[21] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux30( .out( temp4[30] ), .in0( temp3[30] ), .in1( temp3[22] ), .sel( dataB[3] ) ) ;
  Mux_1 B3_Mux31( .out( temp4[31] ), .in0( temp3[31] ), .in1( temp3[23] ), .sel( dataB[3] ) ) ;
  
  Mux_1 B4_Mux0( .out( temp5[0] ), .in0( temp4[0] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux1( .out( temp5[1] ), .in0( temp4[1] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux2( .out( temp5[2] ), .in0( temp4[2] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux3( .out( temp5[3] ), .in0( temp4[3] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux4( .out( temp5[4] ), .in0( temp4[4] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux5( .out( temp5[5] ), .in0( temp4[5] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux6( .out( temp5[6] ), .in0( temp4[6] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux7( .out( temp5[7] ), .in0( temp4[7] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux8( .out( temp5[8] ), .in0( temp4[8] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux9( .out( temp5[9] ), .in0( temp4[9] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux10( .out( temp5[10] ), .in0( temp4[10] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux11( .out( temp5[11] ), .in0( temp4[11] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux12( .out( temp5[12] ), .in0( temp4[12] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux13( .out( temp5[13] ), .in0( temp4[13] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux14( .out( temp5[14] ), .in0( temp4[14] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux15( .out( temp5[15] ), .in0( temp4[15] ), .in1( 1'b0 ), .sel( dataB[4] ) ) ; 
  Mux_1 B4_Mux16( .out( temp5[16] ), .in0( temp4[16] ), .in1( temp4[0] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux17( .out( temp5[17] ), .in0( temp4[17] ), .in1( temp4[1] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux18( .out( temp5[18] ), .in0( temp4[18] ), .in1( temp4[2] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux19( .out( temp5[19] ), .in0( temp4[19] ), .in1( temp4[3] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux20( .out( temp5[20] ), .in0( temp4[20] ), .in1( temp4[4] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux21( .out( temp5[21] ), .in0( temp4[21] ), .in1( temp4[5] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux22( .out( temp5[22] ), .in0( temp4[22] ), .in1( temp4[6] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux23( .out( temp5[23] ), .in0( temp4[23] ), .in1( temp4[7] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux24( .out( temp5[24] ), .in0( temp4[24] ), .in1( temp4[8] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux25( .out( temp5[25] ), .in0( temp4[25] ), .in1( temp4[9] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux26( .out( temp5[26] ), .in0( temp4[26] ), .in1( temp4[10] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux27( .out( temp5[27] ), .in0( temp4[27] ), .in1( temp4[11] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux28( .out( temp5[28] ), .in0( temp4[28] ), .in1( temp4[12] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux29( .out( temp5[29] ), .in0( temp4[29] ), .in1( temp4[13] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux30( .out( temp5[30] ), .in0( temp4[30] ), .in1( temp4[14] ), .sel( dataB[4] ) ) ;
  Mux_1 B4_Mux31( .out( temp5[31] ), .in0( temp4[31] ), .in1( temp4[15] ), .sel( dataB[4] ) ) ;
  
assign dataOut = temp5 ;
endmodule